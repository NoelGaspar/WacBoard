******
* Spice Model
* Item: 1N4148
* Date: 12/07/11
* Revision History: REV A
*==========================================================
* This model was developed by: 
* Central Semiconductor Corp.
* 145 Adams Avenue
* Hauppauge, NY 11788
*
* These models are subject to change without notice.
* Users may not directly or indirectly re-sell or 
* re-distribute this model. This model may not 
* be modified, or altered without the consent of Central Semiconductor Corp. 
*
* For more information on this model contact
* Central Semiconductor Corp. at:
* (631) 435-1110 or Engineering@centralsemi.com
* http://www.centralsemi.com
*==========================================================
******
*SRC=1N4148;1N4148;Diodes;Si;100V  150mA  4.0ns  Central Semi Central Semi
.MODEL 1N4148 D  ( IS=6.2229E-9
+ N=1.9224
+ RS=.33636
+ IKF=42.843E-3
+ CJO=764.38E-15
+ M=.1001
+ VJ=9.9900
+ ISR=11.526E-9
+ NR=4.9950
+ BV=100.14
+ IBV=.25951
+ TT=2.8854E-9 )
******